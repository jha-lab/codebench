module mac_lane_tb();

parameter IL = 4, FL = 16;

logic clk, reset;
logic signed [IL+FL-1:0] i_0, i_1, i_2, i_3, i_4, i_5, i_6, i_7;
logic signed [IL+FL-1:0] i_8, i_9, i_10, i_11, i_12, i_13, i_14, i_15;
logic signed [IL+FL-1:0] w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7;
logic signed [IL+FL-1:0] w_8, w_9, w_10, w_11, w_12, w_13, w_14, w_15;
logic signed [IL+FL-1:0] f;

mac_lane #(.IL(IL), .FL(FL)) mac_lane_0
(
	.clk		(clk),
	.reset		(reset),
	.i_0		(i_0),
	.i_1		(i_1),
	.i_2		(i_2),
	.i_3		(i_3),
	.i_4		(i_4),
	.i_5		(i_5),
	.i_6		(i_6),
	.i_7		(i_7),
	.i_8		(i_8),
	.i_9		(i_9),
	.i_10		(i_10),
	.i_11		(i_11),
	.i_12		(i_12),
	.i_13		(i_13),
	.i_14		(i_14),
	.i_15		(i_15),
	.w_0		(w_0),
	.w_1		(w_1),
	.w_2		(w_2),
	.w_3		(w_3),
	.w_4		(w_4),
	.w_5		(w_5),
	.w_6		(w_6),
	.w_7		(w_7),
	.w_8		(w_8),
	.w_9		(w_9),
	.w_10		(w_10),
	.w_11		(w_11),
	.w_12		(w_12),
	.w_13		(w_13),
	.w_14		(w_14),
	.w_15		(w_15),
	.f		(f)
);

always_ff @(posedge clk) begin
	$display("clk=%b, reset=%b ", clk, reset,
 		 "i_0=%b, i_1=%b, i_2=%b, i_3=%b ", i_0, i_1, i_2, i_3,
		 "i_4=%b, i_5=%b, i_6=%b, i_7=%b ", i_4, i_5, i_6, i_7,
 		 "i_8=%b, i_9=%b, i_10=%b, i_11=%b ", i_8, i_9, i_10, i_11,
 		 "i_12=%b, i_13=%b, i_14=%b, i_15=%b ", i_12, i_13, i_14, i_15,
		 "w_0=%b, w_1=%b, w_2=%b, w_3=%b ", w_0, w_1, w_2, w_3,
 		 "w_4=%b, w_5=%b, w_6=%b, w_7=%b ", w_4, w_5, w_6, w_7,
 		 "w_8=%b, w_9=%b, w_10=%b, w_11=%b ", w_8, w_9, w_10, w_11,
 		 "w_12=%b, w_13=%b, w_14=%b, w_15=%b ", w_12, w_13, w_14, w_15,
 		 "f=%b\n", f);
end


initial begin
	forever begin
		clk = 0;
		#5
		clk = 1;
		#5
		clk = 0;
	end
end

initial begin
	reset = 0;
	i_0 = 20'b0;
	i_1 = 20'b0;
	i_2 = 20'b0;
	i_3 = 20'b0;
	i_4 = 20'b0;
	i_5 = 20'b0;
	i_6 = 20'b0;
	i_7 = 20'b0;
	i_8 = 20'b0;
	i_9 = 20'b0;
	i_10 = 20'b0;
	i_11 = 20'b0;
	i_12 = 20'b0;
	i_13 = 20'b0;
	i_14 = 20'b0;
	i_15 = 20'b0;
	w_0 = 20'b0;
	w_1 = 20'b0;
	w_2 = 20'b0;
	w_3 = 20'b0;
	w_4 = 20'b0;
	w_5 = 20'b0;
	w_6 = 20'b0;
	w_7 = 20'b0;
	w_8 = 20'b0;
	w_9 = 20'b0;
	w_10 = 20'b0;
	w_11 = 20'b0;
	w_12 = 20'b0;
	w_13 = 20'b0;
	w_14 = 20'b0;
	w_15 = 20'b0;
	#50
	reset = 1;
	#50
	reset = 0;
	#100
	i_0 = 20'd0 << 10;
	i_1 = 20'd1 << 10;
	i_2 = 20'd2 << 10;
	i_3 = 20'd3 << 10;
	i_4 = 20'd4 << 10;
	i_5 = 20'd5 << 10;
	i_6 = 20'd6 << 10;
	i_7 = 20'd7 << 10;
	i_8 = 20'd8 << 10;
	i_9 = 20'd9 << 10;
	i_10 = 20'd10 << 10;
	i_11 = 20'd11 << 10;
	i_12 = 20'd12 << 10;
	i_13 = 20'd13 << 10;
	i_14 = 20'd14 << 10;
	i_15 = 20'd15 << 10;
	w_0 = 20'd1 << 10;
	w_1 = 20'd2 << 10;
	w_2 = 20'd3 << 10;
	w_3 = 20'd4 << 10;
	w_4 = 20'd5 << 10;
	w_5 = 20'd6 << 10;
	w_6 = 20'd7 << 10;
	w_7 = 20'd8 << 10;
	w_8 = 20'd9 << 10;
	w_9 = 20'd10 << 10;
	w_10 = 20'd11 << 10;
	w_11 = 20'd12 << 10;
	w_12 = 20'd13 << 10;
	w_13 = 20'd14 << 10;
	w_14 = 20'd15 << 10;
	w_15 = 20'd16 << 10;
	#100
	i_0 = 20'd1 << 10;
	i_1 = 20'd1 << 11;
	i_2 = 20'd1 << 12;
	i_3 = 20'd1 << 13;
	i_4 = 20'd1 << 14;
	i_5 = 20'd1 << 15;
	i_6 = 20'd1 << 10;
	i_7 = 20'd1 << 10;
	i_8 = 20'd0;
	i_9 = 20'd0;
	i_10 = 20'd0;
	i_11 = 20'd0;
	i_12 = 20'd0;
	i_13 = 20'd0;
	i_14 = 20'd0;
	i_15 = 20'd0;
	w_0 = 20'd1 << 10;
	w_1 = 20'd1 << 11;
	w_2 = 20'd1 << 12;
	w_3 = 20'd1 << 13;
	w_4 = 20'd1 << 14;
	w_5 = 20'd1 << 15;
	w_6 = 20'd1 << 10;
	w_7 = 20'd1 << 10;
	w_8 = 20'd1 << 10;
	w_9 = 20'd1 << 10;
	w_10 = 20'd1 << 10;
	w_11 = 20'd1 << 10;
	w_12 = 20'd1 << 10;
	w_13 = 20'd1 << 10;
	w_14 = 20'd1 << 10;
	w_15 = 20'd1 << 10;
	
	#500
	$finish;
	$dumpfile("mac_lane_tb.vcd");
end
endmodule
